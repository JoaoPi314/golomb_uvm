typedef virtual interface_if.mst interface_vif;

class driver extends uvm_driver #(transaction_in);
	`uvm_component_utils(driver) //Sempre tem que ter isso em classes que derivam de uvm_object

	interface_vif vif;
	transaction_in tr;

	function new(string name = "driver", uvm_component parent = null);
		super.new(name, parent);
	endfunction : new


	virtual function void build_phase (uvm_phase phase);
		super.build_phase(phase);
		if(!uvm_config_db#(interface_vif)::get(this, "", "vif", vif))begin
			`uvm_fatal("NOVIF", "failder to get virtual interface")
		end
	endfunction : build_phase

	task run_phase(uvm_phase phase);
		fork
			reset_signals();
			get_and_drive(phase);
		join
	endtask : run_phase

	virtual task reset_signals();
		wait(vif.rstn === 0);
			forever begin
				vif.dt_i    <= '0;
				vif.valid_i <= '0;
				@(posedge vif.rstn);
			end
	endtask : reset_signals


	virtual task get_and_drive(uvm_phase phase);
		wait(vif.rstn === 0);
		@(posedge vif.rstn);
		forever begin
			@(posedge vif.clk);
			seq_item_port.get_next_item(tr);
			$display("dt_i driver= %b", tr.dt_i);
			begin_tr(tr, "req_qdriver");
			@(posedge vif.clk);
			vif.dt_i = tr.dt_i;
			vif.valid_i = '1;
			repeat(2) @(posedge vif.clk);
			vif.valid_i = '0;
			@(negedge vif.busy_o);
			seq_item_port.item_done();
			end_tr(tr);
		end
	endtask : get_and_drive

endclass : driver


